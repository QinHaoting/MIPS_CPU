`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2017/11/02 14:29:33
// Design Name: 
// Module Name: signext
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module signext(
	input wire[15:0] a,
	input wire[1:0] type,
	output wire[31:0] y
    );
	
	// assign y = {{16{a[15]}},a};
	// assign y = {{16{1'b0}}, a};

	// 通过指令的[29:28]判断是否是逻辑运算的立即数扩展
	// “逻辑运算”的立即数0用扩展，而其它立即数用符号位扩展
	assign y = (type == 2'b11) ? {{16{1'b0}}, a} : {{16{a[15]}}, a};
endmodule
